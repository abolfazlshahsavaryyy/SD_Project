-------------------------------------------------------------------------------
--
-- Title       : rotate_register
-- Design      : Shift_Register
-- Author      : abolfazl
-- Company     : google
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\SD_project\Shift_Register\src\rotate_register.vhd
-- Generated   : Sun Aug  3 11:26:59 2025
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {rotate_register} architecture {rotate_register}}



entity rotate_register is
end rotate_register;

--}} End of automatically maintained section

architecture rotate_register of rotate_register is
begin

	 -- enter your statements here --

end rotate_register;
